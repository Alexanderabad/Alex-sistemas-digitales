module led( 
    output z0,
    output z1,
    output z2,
    output z3,
    input a0,
    input b0, 
    input a1,  
    input b1, 
    input a2, 
    input b2, 
    input a3, 
    input b3
);

assign z0 = ~(a0 ^ b0);
assign z1 = ~(a1 ^ b1); 
assign z2 = ~(a2 ^ b2); 
assign z3 = ~(a3 ^ b3);

endmodule